# VerifAI TestGuru
# explain for: axi_adapter.sv
The axi_adapter module implements a simple AXI bus adapter. It supports read and write requests and atomic operations. The module can handle both single and multiple outstanding requests. The module supports cacheline aligned accesses and critical word first accesses. The module also supports wrapping transfers.