# VerifAI TestGuru
# explain for: fpu_wrap.sv
The first part of the code defines the parameters for the floating-point unit. The second part defines the inputs to the FPU and the protocol inversion buffer. The third part translates the inputs.