# VerifAI TestGuru
# explain for: issue_stage.sv
This module implements the issue stage of the RISC-V pipeline. It is responsible for dispatching instructions to the FUs and keeping track of them in a scoreboard like data-structure.