# VerifAI TestGuru
# tests for: instr_realign.sv
```
```