# VerifAI TestGuru
# tests for: load_store_unit.sv
```
```