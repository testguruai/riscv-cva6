# VerifAI TestGuru
# explain for: ex_stage.sv
This module instantiates all functional units residing in the execute stage.