# VerifAI TestGuru
# explain for: cva6.sv
This is the top-level module of the CVA6 core. It instantiates all the modules of the core and connects them together.