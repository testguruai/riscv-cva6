// VerifAI TestGuru
// tests for: compressed_decoder.sv
